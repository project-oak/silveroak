--
-- Copyright 2019 The Project Oak Authors
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--

package and2_package is

  component and2 is
   port(signal a : in bit;
        signal b : bit;
        signal c : out bit);
  end component and2;

end package and2_package;

entity and2 is
 port(signal a : in bit;
      signal b : bit;
      signal c : out bit);
end entity and2;

architecture behavioural of and2 is
begin

 and2_behaviour : process (a) is
   begin
     c <= a and b;
   end process and2_behaviour;

end architecture behavioural;