(****************************************************************************)
(* Copyright 2020 The Project Oak Authors                                   *)
(*                                                                          *)
(* Licensed under the Apache License, Version 2.0 (the "License")           *)
(* you may not use this file except in compliance with the License.         *)
(* You may obtain a copy of the License at                                  *)
(*                                                                          *)
(*     http://www.apache.org/licenses/LICENSE-2.0                           *)
(*                                                                          *)
(* Unless required by applicable law or agreed to in writing, software      *)
(* distributed under the License is distributed on an "AS IS" BASIS,        *)
(* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. *)
(* See the License for the specific language governing permissions and      *)
(* limitations under the License.                                           *)
(****************************************************************************)

From Coq Require Import Arith Eqdep_dec Vector Lia NArith Omega String Ndigits.
From Arrow Require Import Category Arrow.
From Cava Require Import Arrow.ArrowExport BitArithmetic.

From ArrowExamples Require Import Combinators Aes.pkg Aes.sbox.

Import VectorNotations.
Import KappaNotation.
Open Scope kind_scope.

(* module aes_shift_rows (
  input  aes_pkg::ciph_op_e    op_i,
  input  logic [3:0][3:0][7:0] data_i,
  output logic [3:0][3:0][7:0] data_o
); *)
Definition aes_shift_rows
  :  
    <<Bit, Vector (Vector (Vector Bit 8) 4) 4, Unit>> ~> 
      Vector (Vector (Vector Bit 8) 4) 4 :=
  (* // Individually substitute bytes
  import aes_pkg::*;

  // Row 0 is left untouched
  assign data_o[0] = data_i[0];

  // Row 2 does not depend on op_i
  assign data_o[2] = aes_circ_byte_shift(data_i[2], 2'h2);

  // Row 1
  assign data_o[1] = (op_i == CIPH_FWD) ? aes_circ_byte_shift(data_i[1], 2'h3)
                                        : aes_circ_byte_shift(data_i[1], 2'h1);

  // Row 3
  assign data_o[3] = (op_i == CIPH_FWD) ? aes_circ_byte_shift(data_i[3], 2'h1)
                                        : aes_circ_byte_shift(data_i[3], 2'h3); *)
  <[\op_i data_i =>
    let data_o_0 = data_i[#0] in
    let data_o_2 = !aes_circ_byte_shift data_i[#2] (#2) in
    let data_o_1 = 
      if op_i == !CIPH_FWD 
      then !aes_circ_byte_shift data_i[#1] #3
      else !aes_circ_byte_shift data_i[#1] #1
      in
    let data_o_3 = 
      if op_i == !CIPH_FWD 
      then !aes_circ_byte_shift data_i[#3] #1
      else !aes_circ_byte_shift data_i[#3] #3
      in
    data_o_0 :: data_o_1 :: data_o_2 :: data_o_3 :: []
  ]>.

Definition shift_rows_composed :=
  <[\input => 
  let encoded = !aes_shift_rows !CIPH_FWD input in
  let decoded = !aes_shift_rows !CIPH_INV encoded in
  decoded ]>.

Lemma shift_rows_composed_combinational: is_combinational shift_rows_composed.
Proof. simply_combinational. Qed.

(* Notation "# x" := (nat_to_bitvec_sized 8 x) (at level 99). *)

Set Printing Depth 0.

Axiom first_first: forall {x y z w w2} (f: x~>y) (g:y~>z) (h:(Tuple z w)~>w2), first (Arrow:=CircuitArrow) f >>> (first g >>> h) = first (z:=w) (f >>> g) >>> h.
Axiom swap_swap: forall {x y} , swap (A:=CircuitArrow) (x:=x) (y:=y) >>> swap = id.
Axiom first_id: forall {x z w} (f: _ ~> w), first (Arrow:=CircuitArrow) (x:=x)(z:=z) id >>> f = f.
Axiom unassoc_assoc: forall {x y z w} (f: _ ~> w), unassoc (Arrow:=CircuitArrow) (x:=x)(y:=y)(z:=z) >>> assoc >>> f = f.
(* Axiom assoc_unassoc: forall {x z w} , assoc (Arrow:=CircuitArrow) (x:=x)(z:=z) id >>> f = f. *)

Goal exists x, combinational_evaluation shift_rows_composed shift_rows_composed_combinational x = x.
Proof.
  eexists.
  cbv [combinational_evaluation].
  cbv [shift_rows_composed].
  cbv [ClosureConversion.Closure_conversion].
  cbv [ClosureConversion.closure_conversion].
  cbv [ClosureConversion.closure_conversion'].

  (* repeat match goal with
  | |- context [first swap >>> (first swap >>> _)] => rewrite first_first
  end. *)
  repeat rewrite first_first.
  repeat rewrite swap_swap.
  repeat rewrite first_id.

  match goal with
  | |- context [unassoc >>> assoc >>> ?X ] => 
    rewrite (unassoc_assoc X)
  end.

  rewrite (unassoc_assoc _).

  rewrite unassoc_assoc.

  repeat match goal with
  | |- context [first swap >>> (first swap >>> _)] => rewrite first_first
  end.

  
