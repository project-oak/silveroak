package cava is

  component inv is
    port(signal i : in bit;
         signal o : out bit);
  end component inv;

end package cava;